module compuerta_or #(parameter N = 8)(input logic [N-1:0] a,b,
										output logic [N-1:0] or_out );
										
assign or_out = a | b;

endmodule