module compuerta_not #(parameter N = 8)(input logic [N-1:0] a,
													 output logic [N-1:0] not_out );
										
assign not_out = ~a;

endmodule
